`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 09/20/2023 02:24:44 PM
// Design Name: 
// Module Name: ddpls
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module ddpls( input [31:0] a, input  [4:0] b , output  [31:0] o);

assign o = (b == 1)? {a[30:0],a[31]}:
           (b == 2)? {a[29:0],a[31:30]}:
           (b == 3)? {a[28:0],a[31:29]}:
           (b == 4)? {a[27:0],a[31:28]}:
           (b == 5)? {a[26:0],a[31:27]}:
           (b == 6)? {a[25:0],a[31:26]}:
           (b == 7)? {a[24:0],a[31:25]}:
           (b == 8)? {a[23:0],a[31:24]}:
           (b == 9)? {a[22:0],a[31:23]}:
           (b == 10)? {a[21:0],a[31:22]}:
           (b == 11)? {a[20:0],a[31:21]}:
           (b == 12)? {a[19:0],a[31:20]}:
           (b == 13)? {a[18:0],a[31:19]}:
           (b == 14)? {a[17:0],a[31:18]}:
           (b == 15)? {a[16:0],a[31:17]}:
           (b == 16)? {a[15:0],a[31:16]}:
           (b == 17)? {a[14:0],a[31:15]}:
           (b == 18)? {a[13:0],a[31:14]}:
           (b == 19)? {a[12:0],a[31:13]}:
           (b == 20)? {a[11:0],a[31:12]}:
           (b == 21)? {a[10:0],a[31:11]}:
           (b == 22)? {a[9:0],a[31:10]}:
           (b == 23)? {a[8:0],a[31:9]}:
           (b == 24)? {a[7:0],a[31:8]}:
           (b == 25)? {a[6:0],a[31:7]}:
           (b == 26)? {a[5:0],a[31:6]}:
           (b == 27)? {a[4:0],a[31:5]}:
           (b == 28)? {a[3:0],a[31:4]}:
           (b == 29)? {a[2:0],a[31:3]}:
           (b == 30)? {a[1:0],a[31:2]}:
           (b == 31)? {a[0],a[31:1]}:
                      a[31:0];
          

endmodule
